`include "constants.v"
`include "util.v"
module mux1024to1(output [0:`LOG_PORTS_CNT-1]OUT,
				  input [0:9]select,
				  input [0:`TABLE_SIZE-1]TABLE
);

genvar util_genvar;
`MAKE_ARRAY(table_port,TABLE,1000,`LOG_PORTS_CNT,GEN_TABLE_PORT)

assign OUT = (
            select[0:9] == 10'd0 ? table_port[0] :
            select[0:9] == 10'd1 ? table_port[1] :
            select[0:9] == 10'd2 ? table_port[2] :
            select[0:9] == 10'd3 ? table_port[3] :
            select[0:9] == 10'd4 ? table_port[4] :
            select[0:9] == 10'd5 ? table_port[5] :
            select[0:9] == 10'd6 ? table_port[6] :
            select[0:9] == 10'd7 ? table_port[7] :
            select[0:9] == 10'd8 ? table_port[8] :
            select[0:9] == 10'd9 ? table_port[9] :
            select[0:9] == 10'd10 ? table_port[10] :
            select[0:9] == 10'd11 ? table_port[11] :
            select[0:9] == 10'd12 ? table_port[12] :
            select[0:9] == 10'd13 ? table_port[13] :
            select[0:9] == 10'd14 ? table_port[14] :
            select[0:9] == 10'd15 ? table_port[15] :
            select[0:9] == 10'd16 ? table_port[16] :
            select[0:9] == 10'd17 ? table_port[17] :
            select[0:9] == 10'd18 ? table_port[18] :
            select[0:9] == 10'd19 ? table_port[19] :
            select[0:9] == 10'd20 ? table_port[20] :
            select[0:9] == 10'd21 ? table_port[21] :
            select[0:9] == 10'd22 ? table_port[22] :
            select[0:9] == 10'd23 ? table_port[23] :
            select[0:9] == 10'd24 ? table_port[24] :
            select[0:9] == 10'd25 ? table_port[25] :
            select[0:9] == 10'd26 ? table_port[26] :
            select[0:9] == 10'd27 ? table_port[27] :
            select[0:9] == 10'd28 ? table_port[28] :
            select[0:9] == 10'd29 ? table_port[29] :
            select[0:9] == 10'd30 ? table_port[30] :
            select[0:9] == 10'd31 ? table_port[31] :
            select[0:9] == 10'd32 ? table_port[32] :
            select[0:9] == 10'd33 ? table_port[33] :
            select[0:9] == 10'd34 ? table_port[34] :
            select[0:9] == 10'd35 ? table_port[35] :
            select[0:9] == 10'd36 ? table_port[36] :
            select[0:9] == 10'd37 ? table_port[37] :
            select[0:9] == 10'd38 ? table_port[38] :
            select[0:9] == 10'd39 ? table_port[39] :
            select[0:9] == 10'd40 ? table_port[40] :
            select[0:9] == 10'd41 ? table_port[41] :
            select[0:9] == 10'd42 ? table_port[42] :
            select[0:9] == 10'd43 ? table_port[43] :
            select[0:9] == 10'd44 ? table_port[44] :
            select[0:9] == 10'd45 ? table_port[45] :
            select[0:9] == 10'd46 ? table_port[46] :
            select[0:9] == 10'd47 ? table_port[47] :
            select[0:9] == 10'd48 ? table_port[48] :
            select[0:9] == 10'd49 ? table_port[49] :
            select[0:9] == 10'd50 ? table_port[50] :
            select[0:9] == 10'd51 ? table_port[51] :
            select[0:9] == 10'd52 ? table_port[52] :
            select[0:9] == 10'd53 ? table_port[53] :
            select[0:9] == 10'd54 ? table_port[54] :
            select[0:9] == 10'd55 ? table_port[55] :
            select[0:9] == 10'd56 ? table_port[56] :
            select[0:9] == 10'd57 ? table_port[57] :
            select[0:9] == 10'd58 ? table_port[58] :
            select[0:9] == 10'd59 ? table_port[59] :
            select[0:9] == 10'd60 ? table_port[60] :
            select[0:9] == 10'd61 ? table_port[61] :
            select[0:9] == 10'd62 ? table_port[62] :
            select[0:9] == 10'd63 ? table_port[63] :
            select[0:9] == 10'd64 ? table_port[64] :
            select[0:9] == 10'd65 ? table_port[65] :
            select[0:9] == 10'd66 ? table_port[66] :
            select[0:9] == 10'd67 ? table_port[67] :
            select[0:9] == 10'd68 ? table_port[68] :
            select[0:9] == 10'd69 ? table_port[69] :
            select[0:9] == 10'd70 ? table_port[70] :
            select[0:9] == 10'd71 ? table_port[71] :
            select[0:9] == 10'd72 ? table_port[72] :
            select[0:9] == 10'd73 ? table_port[73] :
            select[0:9] == 10'd74 ? table_port[74] :
            select[0:9] == 10'd75 ? table_port[75] :
            select[0:9] == 10'd76 ? table_port[76] :
            select[0:9] == 10'd77 ? table_port[77] :
            select[0:9] == 10'd78 ? table_port[78] :
            select[0:9] == 10'd79 ? table_port[79] :
            select[0:9] == 10'd80 ? table_port[80] :
            select[0:9] == 10'd81 ? table_port[81] :
            select[0:9] == 10'd82 ? table_port[82] :
            select[0:9] == 10'd83 ? table_port[83] :
            select[0:9] == 10'd84 ? table_port[84] :
            select[0:9] == 10'd85 ? table_port[85] :
            select[0:9] == 10'd86 ? table_port[86] :
            select[0:9] == 10'd87 ? table_port[87] :
            select[0:9] == 10'd88 ? table_port[88] :
            select[0:9] == 10'd89 ? table_port[89] :
            select[0:9] == 10'd90 ? table_port[90] :
            select[0:9] == 10'd91 ? table_port[91] :
            select[0:9] == 10'd92 ? table_port[92] :
            select[0:9] == 10'd93 ? table_port[93] :
            select[0:9] == 10'd94 ? table_port[94] :
            select[0:9] == 10'd95 ? table_port[95] :
            select[0:9] == 10'd96 ? table_port[96] :
            select[0:9] == 10'd97 ? table_port[97] :
            select[0:9] == 10'd98 ? table_port[98] :
            select[0:9] == 10'd99 ? table_port[99] :
            select[0:9] == 10'd100 ? table_port[100] :
            select[0:9] == 10'd101 ? table_port[101] :
            select[0:9] == 10'd102 ? table_port[102] :
            select[0:9] == 10'd103 ? table_port[103] :
            select[0:9] == 10'd104 ? table_port[104] :
            select[0:9] == 10'd105 ? table_port[105] :
            select[0:9] == 10'd106 ? table_port[106] :
            select[0:9] == 10'd107 ? table_port[107] :
            select[0:9] == 10'd108 ? table_port[108] :
            select[0:9] == 10'd109 ? table_port[109] :
            select[0:9] == 10'd110 ? table_port[110] :
            select[0:9] == 10'd111 ? table_port[111] :
            select[0:9] == 10'd112 ? table_port[112] :
            select[0:9] == 10'd113 ? table_port[113] :
            select[0:9] == 10'd114 ? table_port[114] :
            select[0:9] == 10'd115 ? table_port[115] :
            select[0:9] == 10'd116 ? table_port[116] :
            select[0:9] == 10'd117 ? table_port[117] :
            select[0:9] == 10'd118 ? table_port[118] :
            select[0:9] == 10'd119 ? table_port[119] :
            select[0:9] == 10'd120 ? table_port[120] :
            select[0:9] == 10'd121 ? table_port[121] :
            select[0:9] == 10'd122 ? table_port[122] :
            select[0:9] == 10'd123 ? table_port[123] :
            select[0:9] == 10'd124 ? table_port[124] :
            select[0:9] == 10'd125 ? table_port[125] :
            select[0:9] == 10'd126 ? table_port[126] :
            select[0:9] == 10'd127 ? table_port[127] :
            select[0:9] == 10'd128 ? table_port[128] :
            select[0:9] == 10'd129 ? table_port[129] :
            select[0:9] == 10'd130 ? table_port[130] :
            select[0:9] == 10'd131 ? table_port[131] :
            select[0:9] == 10'd132 ? table_port[132] :
            select[0:9] == 10'd133 ? table_port[133] :
            select[0:9] == 10'd134 ? table_port[134] :
            select[0:9] == 10'd135 ? table_port[135] :
            select[0:9] == 10'd136 ? table_port[136] :
            select[0:9] == 10'd137 ? table_port[137] :
            select[0:9] == 10'd138 ? table_port[138] :
            select[0:9] == 10'd139 ? table_port[139] :
            select[0:9] == 10'd140 ? table_port[140] :
            select[0:9] == 10'd141 ? table_port[141] :
            select[0:9] == 10'd142 ? table_port[142] :
            select[0:9] == 10'd143 ? table_port[143] :
            select[0:9] == 10'd144 ? table_port[144] :
            select[0:9] == 10'd145 ? table_port[145] :
            select[0:9] == 10'd146 ? table_port[146] :
            select[0:9] == 10'd147 ? table_port[147] :
            select[0:9] == 10'd148 ? table_port[148] :
            select[0:9] == 10'd149 ? table_port[149] :
            select[0:9] == 10'd150 ? table_port[150] :
            select[0:9] == 10'd151 ? table_port[151] :
            select[0:9] == 10'd152 ? table_port[152] :
            select[0:9] == 10'd153 ? table_port[153] :
            select[0:9] == 10'd154 ? table_port[154] :
            select[0:9] == 10'd155 ? table_port[155] :
            select[0:9] == 10'd156 ? table_port[156] :
            select[0:9] == 10'd157 ? table_port[157] :
            select[0:9] == 10'd158 ? table_port[158] :
            select[0:9] == 10'd159 ? table_port[159] :
            select[0:9] == 10'd160 ? table_port[160] :
            select[0:9] == 10'd161 ? table_port[161] :
            select[0:9] == 10'd162 ? table_port[162] :
            select[0:9] == 10'd163 ? table_port[163] :
            select[0:9] == 10'd164 ? table_port[164] :
            select[0:9] == 10'd165 ? table_port[165] :
            select[0:9] == 10'd166 ? table_port[166] :
            select[0:9] == 10'd167 ? table_port[167] :
            select[0:9] == 10'd168 ? table_port[168] :
            select[0:9] == 10'd169 ? table_port[169] :
            select[0:9] == 10'd170 ? table_port[170] :
            select[0:9] == 10'd171 ? table_port[171] :
            select[0:9] == 10'd172 ? table_port[172] :
            select[0:9] == 10'd173 ? table_port[173] :
            select[0:9] == 10'd174 ? table_port[174] :
            select[0:9] == 10'd175 ? table_port[175] :
            select[0:9] == 10'd176 ? table_port[176] :
            select[0:9] == 10'd177 ? table_port[177] :
            select[0:9] == 10'd178 ? table_port[178] :
            select[0:9] == 10'd179 ? table_port[179] :
            select[0:9] == 10'd180 ? table_port[180] :
            select[0:9] == 10'd181 ? table_port[181] :
            select[0:9] == 10'd182 ? table_port[182] :
            select[0:9] == 10'd183 ? table_port[183] :
            select[0:9] == 10'd184 ? table_port[184] :
            select[0:9] == 10'd185 ? table_port[185] :
            select[0:9] == 10'd186 ? table_port[186] :
            select[0:9] == 10'd187 ? table_port[187] :
            select[0:9] == 10'd188 ? table_port[188] :
            select[0:9] == 10'd189 ? table_port[189] :
            select[0:9] == 10'd190 ? table_port[190] :
            select[0:9] == 10'd191 ? table_port[191] :
            select[0:9] == 10'd192 ? table_port[192] :
            select[0:9] == 10'd193 ? table_port[193] :
            select[0:9] == 10'd194 ? table_port[194] :
            select[0:9] == 10'd195 ? table_port[195] :
            select[0:9] == 10'd196 ? table_port[196] :
            select[0:9] == 10'd197 ? table_port[197] :
            select[0:9] == 10'd198 ? table_port[198] :
            select[0:9] == 10'd199 ? table_port[199] :
            select[0:9] == 10'd200 ? table_port[200] :
            select[0:9] == 10'd201 ? table_port[201] :
            select[0:9] == 10'd202 ? table_port[202] :
            select[0:9] == 10'd203 ? table_port[203] :
            select[0:9] == 10'd204 ? table_port[204] :
            select[0:9] == 10'd205 ? table_port[205] :
            select[0:9] == 10'd206 ? table_port[206] :
            select[0:9] == 10'd207 ? table_port[207] :
            select[0:9] == 10'd208 ? table_port[208] :
            select[0:9] == 10'd209 ? table_port[209] :
            select[0:9] == 10'd210 ? table_port[210] :
            select[0:9] == 10'd211 ? table_port[211] :
            select[0:9] == 10'd212 ? table_port[212] :
            select[0:9] == 10'd213 ? table_port[213] :
            select[0:9] == 10'd214 ? table_port[214] :
            select[0:9] == 10'd215 ? table_port[215] :
            select[0:9] == 10'd216 ? table_port[216] :
            select[0:9] == 10'd217 ? table_port[217] :
            select[0:9] == 10'd218 ? table_port[218] :
            select[0:9] == 10'd219 ? table_port[219] :
            select[0:9] == 10'd220 ? table_port[220] :
            select[0:9] == 10'd221 ? table_port[221] :
            select[0:9] == 10'd222 ? table_port[222] :
            select[0:9] == 10'd223 ? table_port[223] :
            select[0:9] == 10'd224 ? table_port[224] :
            select[0:9] == 10'd225 ? table_port[225] :
            select[0:9] == 10'd226 ? table_port[226] :
            select[0:9] == 10'd227 ? table_port[227] :
            select[0:9] == 10'd228 ? table_port[228] :
            select[0:9] == 10'd229 ? table_port[229] :
            select[0:9] == 10'd230 ? table_port[230] :
            select[0:9] == 10'd231 ? table_port[231] :
            select[0:9] == 10'd232 ? table_port[232] :
            select[0:9] == 10'd233 ? table_port[233] :
            select[0:9] == 10'd234 ? table_port[234] :
            select[0:9] == 10'd235 ? table_port[235] :
            select[0:9] == 10'd236 ? table_port[236] :
            select[0:9] == 10'd237 ? table_port[237] :
            select[0:9] == 10'd238 ? table_port[238] :
            select[0:9] == 10'd239 ? table_port[239] :
            select[0:9] == 10'd240 ? table_port[240] :
            select[0:9] == 10'd241 ? table_port[241] :
            select[0:9] == 10'd242 ? table_port[242] :
            select[0:9] == 10'd243 ? table_port[243] :
            select[0:9] == 10'd244 ? table_port[244] :
            select[0:9] == 10'd245 ? table_port[245] :
            select[0:9] == 10'd246 ? table_port[246] :
            select[0:9] == 10'd247 ? table_port[247] :
            select[0:9] == 10'd248 ? table_port[248] :
            select[0:9] == 10'd249 ? table_port[249] :
            select[0:9] == 10'd250 ? table_port[250] :
            select[0:9] == 10'd251 ? table_port[251] :
            select[0:9] == 10'd252 ? table_port[252] :
            select[0:9] == 10'd253 ? table_port[253] :
            select[0:9] == 10'd254 ? table_port[254] :
            select[0:9] == 10'd255 ? table_port[255] :
            select[0:9] == 10'd256 ? table_port[256] :
            select[0:9] == 10'd257 ? table_port[257] :
            select[0:9] == 10'd258 ? table_port[258] :
            select[0:9] == 10'd259 ? table_port[259] :
            select[0:9] == 10'd260 ? table_port[260] :
            select[0:9] == 10'd261 ? table_port[261] :
            select[0:9] == 10'd262 ? table_port[262] :
            select[0:9] == 10'd263 ? table_port[263] :
            select[0:9] == 10'd264 ? table_port[264] :
            select[0:9] == 10'd265 ? table_port[265] :
            select[0:9] == 10'd266 ? table_port[266] :
            select[0:9] == 10'd267 ? table_port[267] :
            select[0:9] == 10'd268 ? table_port[268] :
            select[0:9] == 10'd269 ? table_port[269] :
            select[0:9] == 10'd270 ? table_port[270] :
            select[0:9] == 10'd271 ? table_port[271] :
            select[0:9] == 10'd272 ? table_port[272] :
            select[0:9] == 10'd273 ? table_port[273] :
            select[0:9] == 10'd274 ? table_port[274] :
            select[0:9] == 10'd275 ? table_port[275] :
            select[0:9] == 10'd276 ? table_port[276] :
            select[0:9] == 10'd277 ? table_port[277] :
            select[0:9] == 10'd278 ? table_port[278] :
            select[0:9] == 10'd279 ? table_port[279] :
            select[0:9] == 10'd280 ? table_port[280] :
            select[0:9] == 10'd281 ? table_port[281] :
            select[0:9] == 10'd282 ? table_port[282] :
            select[0:9] == 10'd283 ? table_port[283] :
            select[0:9] == 10'd284 ? table_port[284] :
            select[0:9] == 10'd285 ? table_port[285] :
            select[0:9] == 10'd286 ? table_port[286] :
            select[0:9] == 10'd287 ? table_port[287] :
            select[0:9] == 10'd288 ? table_port[288] :
            select[0:9] == 10'd289 ? table_port[289] :
            select[0:9] == 10'd290 ? table_port[290] :
            select[0:9] == 10'd291 ? table_port[291] :
            select[0:9] == 10'd292 ? table_port[292] :
            select[0:9] == 10'd293 ? table_port[293] :
            select[0:9] == 10'd294 ? table_port[294] :
            select[0:9] == 10'd295 ? table_port[295] :
            select[0:9] == 10'd296 ? table_port[296] :
            select[0:9] == 10'd297 ? table_port[297] :
            select[0:9] == 10'd298 ? table_port[298] :
            select[0:9] == 10'd299 ? table_port[299] :
            select[0:9] == 10'd300 ? table_port[300] :
            select[0:9] == 10'd301 ? table_port[301] :
            select[0:9] == 10'd302 ? table_port[302] :
            select[0:9] == 10'd303 ? table_port[303] :
            select[0:9] == 10'd304 ? table_port[304] :
            select[0:9] == 10'd305 ? table_port[305] :
            select[0:9] == 10'd306 ? table_port[306] :
            select[0:9] == 10'd307 ? table_port[307] :
            select[0:9] == 10'd308 ? table_port[308] :
            select[0:9] == 10'd309 ? table_port[309] :
            select[0:9] == 10'd310 ? table_port[310] :
            select[0:9] == 10'd311 ? table_port[311] :
            select[0:9] == 10'd312 ? table_port[312] :
            select[0:9] == 10'd313 ? table_port[313] :
            select[0:9] == 10'd314 ? table_port[314] :
            select[0:9] == 10'd315 ? table_port[315] :
            select[0:9] == 10'd316 ? table_port[316] :
            select[0:9] == 10'd317 ? table_port[317] :
            select[0:9] == 10'd318 ? table_port[318] :
            select[0:9] == 10'd319 ? table_port[319] :
            select[0:9] == 10'd320 ? table_port[320] :
            select[0:9] == 10'd321 ? table_port[321] :
            select[0:9] == 10'd322 ? table_port[322] :
            select[0:9] == 10'd323 ? table_port[323] :
            select[0:9] == 10'd324 ? table_port[324] :
            select[0:9] == 10'd325 ? table_port[325] :
            select[0:9] == 10'd326 ? table_port[326] :
            select[0:9] == 10'd327 ? table_port[327] :
            select[0:9] == 10'd328 ? table_port[328] :
            select[0:9] == 10'd329 ? table_port[329] :
            select[0:9] == 10'd330 ? table_port[330] :
            select[0:9] == 10'd331 ? table_port[331] :
            select[0:9] == 10'd332 ? table_port[332] :
            select[0:9] == 10'd333 ? table_port[333] :
            select[0:9] == 10'd334 ? table_port[334] :
            select[0:9] == 10'd335 ? table_port[335] :
            select[0:9] == 10'd336 ? table_port[336] :
            select[0:9] == 10'd337 ? table_port[337] :
            select[0:9] == 10'd338 ? table_port[338] :
            select[0:9] == 10'd339 ? table_port[339] :
            select[0:9] == 10'd340 ? table_port[340] :
            select[0:9] == 10'd341 ? table_port[341] :
            select[0:9] == 10'd342 ? table_port[342] :
            select[0:9] == 10'd343 ? table_port[343] :
            select[0:9] == 10'd344 ? table_port[344] :
            select[0:9] == 10'd345 ? table_port[345] :
            select[0:9] == 10'd346 ? table_port[346] :
            select[0:9] == 10'd347 ? table_port[347] :
            select[0:9] == 10'd348 ? table_port[348] :
            select[0:9] == 10'd349 ? table_port[349] :
            select[0:9] == 10'd350 ? table_port[350] :
            select[0:9] == 10'd351 ? table_port[351] :
            select[0:9] == 10'd352 ? table_port[352] :
            select[0:9] == 10'd353 ? table_port[353] :
            select[0:9] == 10'd354 ? table_port[354] :
            select[0:9] == 10'd355 ? table_port[355] :
            select[0:9] == 10'd356 ? table_port[356] :
            select[0:9] == 10'd357 ? table_port[357] :
            select[0:9] == 10'd358 ? table_port[358] :
            select[0:9] == 10'd359 ? table_port[359] :
            select[0:9] == 10'd360 ? table_port[360] :
            select[0:9] == 10'd361 ? table_port[361] :
            select[0:9] == 10'd362 ? table_port[362] :
            select[0:9] == 10'd363 ? table_port[363] :
            select[0:9] == 10'd364 ? table_port[364] :
            select[0:9] == 10'd365 ? table_port[365] :
            select[0:9] == 10'd366 ? table_port[366] :
            select[0:9] == 10'd367 ? table_port[367] :
            select[0:9] == 10'd368 ? table_port[368] :
            select[0:9] == 10'd369 ? table_port[369] :
            select[0:9] == 10'd370 ? table_port[370] :
            select[0:9] == 10'd371 ? table_port[371] :
            select[0:9] == 10'd372 ? table_port[372] :
            select[0:9] == 10'd373 ? table_port[373] :
            select[0:9] == 10'd374 ? table_port[374] :
            select[0:9] == 10'd375 ? table_port[375] :
            select[0:9] == 10'd376 ? table_port[376] :
            select[0:9] == 10'd377 ? table_port[377] :
            select[0:9] == 10'd378 ? table_port[378] :
            select[0:9] == 10'd379 ? table_port[379] :
            select[0:9] == 10'd380 ? table_port[380] :
            select[0:9] == 10'd381 ? table_port[381] :
            select[0:9] == 10'd382 ? table_port[382] :
            select[0:9] == 10'd383 ? table_port[383] :
            select[0:9] == 10'd384 ? table_port[384] :
            select[0:9] == 10'd385 ? table_port[385] :
            select[0:9] == 10'd386 ? table_port[386] :
            select[0:9] == 10'd387 ? table_port[387] :
            select[0:9] == 10'd388 ? table_port[388] :
            select[0:9] == 10'd389 ? table_port[389] :
            select[0:9] == 10'd390 ? table_port[390] :
            select[0:9] == 10'd391 ? table_port[391] :
            select[0:9] == 10'd392 ? table_port[392] :
            select[0:9] == 10'd393 ? table_port[393] :
            select[0:9] == 10'd394 ? table_port[394] :
            select[0:9] == 10'd395 ? table_port[395] :
            select[0:9] == 10'd396 ? table_port[396] :
            select[0:9] == 10'd397 ? table_port[397] :
            select[0:9] == 10'd398 ? table_port[398] :
            select[0:9] == 10'd399 ? table_port[399] :
            select[0:9] == 10'd400 ? table_port[400] :
            select[0:9] == 10'd401 ? table_port[401] :
            select[0:9] == 10'd402 ? table_port[402] :
            select[0:9] == 10'd403 ? table_port[403] :
            select[0:9] == 10'd404 ? table_port[404] :
            select[0:9] == 10'd405 ? table_port[405] :
            select[0:9] == 10'd406 ? table_port[406] :
            select[0:9] == 10'd407 ? table_port[407] :
            select[0:9] == 10'd408 ? table_port[408] :
            select[0:9] == 10'd409 ? table_port[409] :
            select[0:9] == 10'd410 ? table_port[410] :
            select[0:9] == 10'd411 ? table_port[411] :
            select[0:9] == 10'd412 ? table_port[412] :
            select[0:9] == 10'd413 ? table_port[413] :
            select[0:9] == 10'd414 ? table_port[414] :
            select[0:9] == 10'd415 ? table_port[415] :
            select[0:9] == 10'd416 ? table_port[416] :
            select[0:9] == 10'd417 ? table_port[417] :
            select[0:9] == 10'd418 ? table_port[418] :
            select[0:9] == 10'd419 ? table_port[419] :
            select[0:9] == 10'd420 ? table_port[420] :
            select[0:9] == 10'd421 ? table_port[421] :
            select[0:9] == 10'd422 ? table_port[422] :
            select[0:9] == 10'd423 ? table_port[423] :
            select[0:9] == 10'd424 ? table_port[424] :
            select[0:9] == 10'd425 ? table_port[425] :
            select[0:9] == 10'd426 ? table_port[426] :
            select[0:9] == 10'd427 ? table_port[427] :
            select[0:9] == 10'd428 ? table_port[428] :
            select[0:9] == 10'd429 ? table_port[429] :
            select[0:9] == 10'd430 ? table_port[430] :
            select[0:9] == 10'd431 ? table_port[431] :
            select[0:9] == 10'd432 ? table_port[432] :
            select[0:9] == 10'd433 ? table_port[433] :
            select[0:9] == 10'd434 ? table_port[434] :
            select[0:9] == 10'd435 ? table_port[435] :
            select[0:9] == 10'd436 ? table_port[436] :
            select[0:9] == 10'd437 ? table_port[437] :
            select[0:9] == 10'd438 ? table_port[438] :
            select[0:9] == 10'd439 ? table_port[439] :
            select[0:9] == 10'd440 ? table_port[440] :
            select[0:9] == 10'd441 ? table_port[441] :
            select[0:9] == 10'd442 ? table_port[442] :
            select[0:9] == 10'd443 ? table_port[443] :
            select[0:9] == 10'd444 ? table_port[444] :
            select[0:9] == 10'd445 ? table_port[445] :
            select[0:9] == 10'd446 ? table_port[446] :
            select[0:9] == 10'd447 ? table_port[447] :
            select[0:9] == 10'd448 ? table_port[448] :
            select[0:9] == 10'd449 ? table_port[449] :
            select[0:9] == 10'd450 ? table_port[450] :
            select[0:9] == 10'd451 ? table_port[451] :
            select[0:9] == 10'd452 ? table_port[452] :
            select[0:9] == 10'd453 ? table_port[453] :
            select[0:9] == 10'd454 ? table_port[454] :
            select[0:9] == 10'd455 ? table_port[455] :
            select[0:9] == 10'd456 ? table_port[456] :
            select[0:9] == 10'd457 ? table_port[457] :
            select[0:9] == 10'd458 ? table_port[458] :
            select[0:9] == 10'd459 ? table_port[459] :
            select[0:9] == 10'd460 ? table_port[460] :
            select[0:9] == 10'd461 ? table_port[461] :
            select[0:9] == 10'd462 ? table_port[462] :
            select[0:9] == 10'd463 ? table_port[463] :
            select[0:9] == 10'd464 ? table_port[464] :
            select[0:9] == 10'd465 ? table_port[465] :
            select[0:9] == 10'd466 ? table_port[466] :
            select[0:9] == 10'd467 ? table_port[467] :
            select[0:9] == 10'd468 ? table_port[468] :
            select[0:9] == 10'd469 ? table_port[469] :
            select[0:9] == 10'd470 ? table_port[470] :
            select[0:9] == 10'd471 ? table_port[471] :
            select[0:9] == 10'd472 ? table_port[472] :
            select[0:9] == 10'd473 ? table_port[473] :
            select[0:9] == 10'd474 ? table_port[474] :
            select[0:9] == 10'd475 ? table_port[475] :
            select[0:9] == 10'd476 ? table_port[476] :
            select[0:9] == 10'd477 ? table_port[477] :
            select[0:9] == 10'd478 ? table_port[478] :
            select[0:9] == 10'd479 ? table_port[479] :
            select[0:9] == 10'd480 ? table_port[480] :
            select[0:9] == 10'd481 ? table_port[481] :
            select[0:9] == 10'd482 ? table_port[482] :
            select[0:9] == 10'd483 ? table_port[483] :
            select[0:9] == 10'd484 ? table_port[484] :
            select[0:9] == 10'd485 ? table_port[485] :
            select[0:9] == 10'd486 ? table_port[486] :
            select[0:9] == 10'd487 ? table_port[487] :
            select[0:9] == 10'd488 ? table_port[488] :
            select[0:9] == 10'd489 ? table_port[489] :
            select[0:9] == 10'd490 ? table_port[490] :
            select[0:9] == 10'd491 ? table_port[491] :
            select[0:9] == 10'd492 ? table_port[492] :
            select[0:9] == 10'd493 ? table_port[493] :
            select[0:9] == 10'd494 ? table_port[494] :
            select[0:9] == 10'd495 ? table_port[495] :
            select[0:9] == 10'd496 ? table_port[496] :
            select[0:9] == 10'd497 ? table_port[497] :
            select[0:9] == 10'd498 ? table_port[498] :
            select[0:9] == 10'd499 ? table_port[499] :
            select[0:9] == 10'd500 ? table_port[500] :
            select[0:9] == 10'd501 ? table_port[501] :
            select[0:9] == 10'd502 ? table_port[502] :
            select[0:9] == 10'd503 ? table_port[503] :
            select[0:9] == 10'd504 ? table_port[504] :
            select[0:9] == 10'd505 ? table_port[505] :
            select[0:9] == 10'd506 ? table_port[506] :
            select[0:9] == 10'd507 ? table_port[507] :
            select[0:9] == 10'd508 ? table_port[508] :
            select[0:9] == 10'd509 ? table_port[509] :
            select[0:9] == 10'd510 ? table_port[510] :
            select[0:9] == 10'd511 ? table_port[511] :
            select[0:9] == 10'd512 ? table_port[512] :
            select[0:9] == 10'd513 ? table_port[513] :
            select[0:9] == 10'd514 ? table_port[514] :
            select[0:9] == 10'd515 ? table_port[515] :
            select[0:9] == 10'd516 ? table_port[516] :
            select[0:9] == 10'd517 ? table_port[517] :
            select[0:9] == 10'd518 ? table_port[518] :
            select[0:9] == 10'd519 ? table_port[519] :
            select[0:9] == 10'd520 ? table_port[520] :
            select[0:9] == 10'd521 ? table_port[521] :
            select[0:9] == 10'd522 ? table_port[522] :
            select[0:9] == 10'd523 ? table_port[523] :
            select[0:9] == 10'd524 ? table_port[524] :
            select[0:9] == 10'd525 ? table_port[525] :
            select[0:9] == 10'd526 ? table_port[526] :
            select[0:9] == 10'd527 ? table_port[527] :
            select[0:9] == 10'd528 ? table_port[528] :
            select[0:9] == 10'd529 ? table_port[529] :
            select[0:9] == 10'd530 ? table_port[530] :
            select[0:9] == 10'd531 ? table_port[531] :
            select[0:9] == 10'd532 ? table_port[532] :
            select[0:9] == 10'd533 ? table_port[533] :
            select[0:9] == 10'd534 ? table_port[534] :
            select[0:9] == 10'd535 ? table_port[535] :
            select[0:9] == 10'd536 ? table_port[536] :
            select[0:9] == 10'd537 ? table_port[537] :
            select[0:9] == 10'd538 ? table_port[538] :
            select[0:9] == 10'd539 ? table_port[539] :
            select[0:9] == 10'd540 ? table_port[540] :
            select[0:9] == 10'd541 ? table_port[541] :
            select[0:9] == 10'd542 ? table_port[542] :
            select[0:9] == 10'd543 ? table_port[543] :
            select[0:9] == 10'd544 ? table_port[544] :
            select[0:9] == 10'd545 ? table_port[545] :
            select[0:9] == 10'd546 ? table_port[546] :
            select[0:9] == 10'd547 ? table_port[547] :
            select[0:9] == 10'd548 ? table_port[548] :
            select[0:9] == 10'd549 ? table_port[549] :
            select[0:9] == 10'd550 ? table_port[550] :
            select[0:9] == 10'd551 ? table_port[551] :
            select[0:9] == 10'd552 ? table_port[552] :
            select[0:9] == 10'd553 ? table_port[553] :
            select[0:9] == 10'd554 ? table_port[554] :
            select[0:9] == 10'd555 ? table_port[555] :
            select[0:9] == 10'd556 ? table_port[556] :
            select[0:9] == 10'd557 ? table_port[557] :
            select[0:9] == 10'd558 ? table_port[558] :
            select[0:9] == 10'd559 ? table_port[559] :
            select[0:9] == 10'd560 ? table_port[560] :
            select[0:9] == 10'd561 ? table_port[561] :
            select[0:9] == 10'd562 ? table_port[562] :
            select[0:9] == 10'd563 ? table_port[563] :
            select[0:9] == 10'd564 ? table_port[564] :
            select[0:9] == 10'd565 ? table_port[565] :
            select[0:9] == 10'd566 ? table_port[566] :
            select[0:9] == 10'd567 ? table_port[567] :
            select[0:9] == 10'd568 ? table_port[568] :
            select[0:9] == 10'd569 ? table_port[569] :
            select[0:9] == 10'd570 ? table_port[570] :
            select[0:9] == 10'd571 ? table_port[571] :
            select[0:9] == 10'd572 ? table_port[572] :
            select[0:9] == 10'd573 ? table_port[573] :
            select[0:9] == 10'd574 ? table_port[574] :
            select[0:9] == 10'd575 ? table_port[575] :
            select[0:9] == 10'd576 ? table_port[576] :
            select[0:9] == 10'd577 ? table_port[577] :
            select[0:9] == 10'd578 ? table_port[578] :
            select[0:9] == 10'd579 ? table_port[579] :
            select[0:9] == 10'd580 ? table_port[580] :
            select[0:9] == 10'd581 ? table_port[581] :
            select[0:9] == 10'd582 ? table_port[582] :
            select[0:9] == 10'd583 ? table_port[583] :
            select[0:9] == 10'd584 ? table_port[584] :
            select[0:9] == 10'd585 ? table_port[585] :
            select[0:9] == 10'd586 ? table_port[586] :
            select[0:9] == 10'd587 ? table_port[587] :
            select[0:9] == 10'd588 ? table_port[588] :
            select[0:9] == 10'd589 ? table_port[589] :
            select[0:9] == 10'd590 ? table_port[590] :
            select[0:9] == 10'd591 ? table_port[591] :
            select[0:9] == 10'd592 ? table_port[592] :
            select[0:9] == 10'd593 ? table_port[593] :
            select[0:9] == 10'd594 ? table_port[594] :
            select[0:9] == 10'd595 ? table_port[595] :
            select[0:9] == 10'd596 ? table_port[596] :
            select[0:9] == 10'd597 ? table_port[597] :
            select[0:9] == 10'd598 ? table_port[598] :
            select[0:9] == 10'd599 ? table_port[599] :
            select[0:9] == 10'd600 ? table_port[600] :
            select[0:9] == 10'd601 ? table_port[601] :
            select[0:9] == 10'd602 ? table_port[602] :
            select[0:9] == 10'd603 ? table_port[603] :
            select[0:9] == 10'd604 ? table_port[604] :
            select[0:9] == 10'd605 ? table_port[605] :
            select[0:9] == 10'd606 ? table_port[606] :
            select[0:9] == 10'd607 ? table_port[607] :
            select[0:9] == 10'd608 ? table_port[608] :
            select[0:9] == 10'd609 ? table_port[609] :
            select[0:9] == 10'd610 ? table_port[610] :
            select[0:9] == 10'd611 ? table_port[611] :
            select[0:9] == 10'd612 ? table_port[612] :
            select[0:9] == 10'd613 ? table_port[613] :
            select[0:9] == 10'd614 ? table_port[614] :
            select[0:9] == 10'd615 ? table_port[615] :
            select[0:9] == 10'd616 ? table_port[616] :
            select[0:9] == 10'd617 ? table_port[617] :
            select[0:9] == 10'd618 ? table_port[618] :
            select[0:9] == 10'd619 ? table_port[619] :
            select[0:9] == 10'd620 ? table_port[620] :
            select[0:9] == 10'd621 ? table_port[621] :
            select[0:9] == 10'd622 ? table_port[622] :
            select[0:9] == 10'd623 ? table_port[623] :
            select[0:9] == 10'd624 ? table_port[624] :
            select[0:9] == 10'd625 ? table_port[625] :
            select[0:9] == 10'd626 ? table_port[626] :
            select[0:9] == 10'd627 ? table_port[627] :
            select[0:9] == 10'd628 ? table_port[628] :
            select[0:9] == 10'd629 ? table_port[629] :
            select[0:9] == 10'd630 ? table_port[630] :
            select[0:9] == 10'd631 ? table_port[631] :
            select[0:9] == 10'd632 ? table_port[632] :
            select[0:9] == 10'd633 ? table_port[633] :
            select[0:9] == 10'd634 ? table_port[634] :
            select[0:9] == 10'd635 ? table_port[635] :
            select[0:9] == 10'd636 ? table_port[636] :
            select[0:9] == 10'd637 ? table_port[637] :
            select[0:9] == 10'd638 ? table_port[638] :
            select[0:9] == 10'd639 ? table_port[639] :
            select[0:9] == 10'd640 ? table_port[640] :
            select[0:9] == 10'd641 ? table_port[641] :
            select[0:9] == 10'd642 ? table_port[642] :
            select[0:9] == 10'd643 ? table_port[643] :
            select[0:9] == 10'd644 ? table_port[644] :
            select[0:9] == 10'd645 ? table_port[645] :
            select[0:9] == 10'd646 ? table_port[646] :
            select[0:9] == 10'd647 ? table_port[647] :
            select[0:9] == 10'd648 ? table_port[648] :
            select[0:9] == 10'd649 ? table_port[649] :
            select[0:9] == 10'd650 ? table_port[650] :
            select[0:9] == 10'd651 ? table_port[651] :
            select[0:9] == 10'd652 ? table_port[652] :
            select[0:9] == 10'd653 ? table_port[653] :
            select[0:9] == 10'd654 ? table_port[654] :
            select[0:9] == 10'd655 ? table_port[655] :
            select[0:9] == 10'd656 ? table_port[656] :
            select[0:9] == 10'd657 ? table_port[657] :
            select[0:9] == 10'd658 ? table_port[658] :
            select[0:9] == 10'd659 ? table_port[659] :
            select[0:9] == 10'd660 ? table_port[660] :
            select[0:9] == 10'd661 ? table_port[661] :
            select[0:9] == 10'd662 ? table_port[662] :
            select[0:9] == 10'd663 ? table_port[663] :
            select[0:9] == 10'd664 ? table_port[664] :
            select[0:9] == 10'd665 ? table_port[665] :
            select[0:9] == 10'd666 ? table_port[666] :
            select[0:9] == 10'd667 ? table_port[667] :
            select[0:9] == 10'd668 ? table_port[668] :
            select[0:9] == 10'd669 ? table_port[669] :
            select[0:9] == 10'd670 ? table_port[670] :
            select[0:9] == 10'd671 ? table_port[671] :
            select[0:9] == 10'd672 ? table_port[672] :
            select[0:9] == 10'd673 ? table_port[673] :
            select[0:9] == 10'd674 ? table_port[674] :
            select[0:9] == 10'd675 ? table_port[675] :
            select[0:9] == 10'd676 ? table_port[676] :
            select[0:9] == 10'd677 ? table_port[677] :
            select[0:9] == 10'd678 ? table_port[678] :
            select[0:9] == 10'd679 ? table_port[679] :
            select[0:9] == 10'd680 ? table_port[680] :
            select[0:9] == 10'd681 ? table_port[681] :
            select[0:9] == 10'd682 ? table_port[682] :
            select[0:9] == 10'd683 ? table_port[683] :
            select[0:9] == 10'd684 ? table_port[684] :
            select[0:9] == 10'd685 ? table_port[685] :
            select[0:9] == 10'd686 ? table_port[686] :
            select[0:9] == 10'd687 ? table_port[687] :
            select[0:9] == 10'd688 ? table_port[688] :
            select[0:9] == 10'd689 ? table_port[689] :
            select[0:9] == 10'd690 ? table_port[690] :
            select[0:9] == 10'd691 ? table_port[691] :
            select[0:9] == 10'd692 ? table_port[692] :
            select[0:9] == 10'd693 ? table_port[693] :
            select[0:9] == 10'd694 ? table_port[694] :
            select[0:9] == 10'd695 ? table_port[695] :
            select[0:9] == 10'd696 ? table_port[696] :
            select[0:9] == 10'd697 ? table_port[697] :
            select[0:9] == 10'd698 ? table_port[698] :
            select[0:9] == 10'd699 ? table_port[699] :
            select[0:9] == 10'd700 ? table_port[700] :
            select[0:9] == 10'd701 ? table_port[701] :
            select[0:9] == 10'd702 ? table_port[702] :
            select[0:9] == 10'd703 ? table_port[703] :
            select[0:9] == 10'd704 ? table_port[704] :
            select[0:9] == 10'd705 ? table_port[705] :
            select[0:9] == 10'd706 ? table_port[706] :
            select[0:9] == 10'd707 ? table_port[707] :
            select[0:9] == 10'd708 ? table_port[708] :
            select[0:9] == 10'd709 ? table_port[709] :
            select[0:9] == 10'd710 ? table_port[710] :
            select[0:9] == 10'd711 ? table_port[711] :
            select[0:9] == 10'd712 ? table_port[712] :
            select[0:9] == 10'd713 ? table_port[713] :
            select[0:9] == 10'd714 ? table_port[714] :
            select[0:9] == 10'd715 ? table_port[715] :
            select[0:9] == 10'd716 ? table_port[716] :
            select[0:9] == 10'd717 ? table_port[717] :
            select[0:9] == 10'd718 ? table_port[718] :
            select[0:9] == 10'd719 ? table_port[719] :
            select[0:9] == 10'd720 ? table_port[720] :
            select[0:9] == 10'd721 ? table_port[721] :
            select[0:9] == 10'd722 ? table_port[722] :
            select[0:9] == 10'd723 ? table_port[723] :
            select[0:9] == 10'd724 ? table_port[724] :
            select[0:9] == 10'd725 ? table_port[725] :
            select[0:9] == 10'd726 ? table_port[726] :
            select[0:9] == 10'd727 ? table_port[727] :
            select[0:9] == 10'd728 ? table_port[728] :
            select[0:9] == 10'd729 ? table_port[729] :
            select[0:9] == 10'd730 ? table_port[730] :
            select[0:9] == 10'd731 ? table_port[731] :
            select[0:9] == 10'd732 ? table_port[732] :
            select[0:9] == 10'd733 ? table_port[733] :
            select[0:9] == 10'd734 ? table_port[734] :
            select[0:9] == 10'd735 ? table_port[735] :
            select[0:9] == 10'd736 ? table_port[736] :
            select[0:9] == 10'd737 ? table_port[737] :
            select[0:9] == 10'd738 ? table_port[738] :
            select[0:9] == 10'd739 ? table_port[739] :
            select[0:9] == 10'd740 ? table_port[740] :
            select[0:9] == 10'd741 ? table_port[741] :
            select[0:9] == 10'd742 ? table_port[742] :
            select[0:9] == 10'd743 ? table_port[743] :
            select[0:9] == 10'd744 ? table_port[744] :
            select[0:9] == 10'd745 ? table_port[745] :
            select[0:9] == 10'd746 ? table_port[746] :
            select[0:9] == 10'd747 ? table_port[747] :
            select[0:9] == 10'd748 ? table_port[748] :
            select[0:9] == 10'd749 ? table_port[749] :
            select[0:9] == 10'd750 ? table_port[750] :
            select[0:9] == 10'd751 ? table_port[751] :
            select[0:9] == 10'd752 ? table_port[752] :
            select[0:9] == 10'd753 ? table_port[753] :
            select[0:9] == 10'd754 ? table_port[754] :
            select[0:9] == 10'd755 ? table_port[755] :
            select[0:9] == 10'd756 ? table_port[756] :
            select[0:9] == 10'd757 ? table_port[757] :
            select[0:9] == 10'd758 ? table_port[758] :
            select[0:9] == 10'd759 ? table_port[759] :
            select[0:9] == 10'd760 ? table_port[760] :
            select[0:9] == 10'd761 ? table_port[761] :
            select[0:9] == 10'd762 ? table_port[762] :
            select[0:9] == 10'd763 ? table_port[763] :
            select[0:9] == 10'd764 ? table_port[764] :
            select[0:9] == 10'd765 ? table_port[765] :
            select[0:9] == 10'd766 ? table_port[766] :
            select[0:9] == 10'd767 ? table_port[767] :
            select[0:9] == 10'd768 ? table_port[768] :
            select[0:9] == 10'd769 ? table_port[769] :
            select[0:9] == 10'd770 ? table_port[770] :
            select[0:9] == 10'd771 ? table_port[771] :
            select[0:9] == 10'd772 ? table_port[772] :
            select[0:9] == 10'd773 ? table_port[773] :
            select[0:9] == 10'd774 ? table_port[774] :
            select[0:9] == 10'd775 ? table_port[775] :
            select[0:9] == 10'd776 ? table_port[776] :
            select[0:9] == 10'd777 ? table_port[777] :
            select[0:9] == 10'd778 ? table_port[778] :
            select[0:9] == 10'd779 ? table_port[779] :
            select[0:9] == 10'd780 ? table_port[780] :
            select[0:9] == 10'd781 ? table_port[781] :
            select[0:9] == 10'd782 ? table_port[782] :
            select[0:9] == 10'd783 ? table_port[783] :
            select[0:9] == 10'd784 ? table_port[784] :
            select[0:9] == 10'd785 ? table_port[785] :
            select[0:9] == 10'd786 ? table_port[786] :
            select[0:9] == 10'd787 ? table_port[787] :
            select[0:9] == 10'd788 ? table_port[788] :
            select[0:9] == 10'd789 ? table_port[789] :
            select[0:9] == 10'd790 ? table_port[790] :
            select[0:9] == 10'd791 ? table_port[791] :
            select[0:9] == 10'd792 ? table_port[792] :
            select[0:9] == 10'd793 ? table_port[793] :
            select[0:9] == 10'd794 ? table_port[794] :
            select[0:9] == 10'd795 ? table_port[795] :
            select[0:9] == 10'd796 ? table_port[796] :
            select[0:9] == 10'd797 ? table_port[797] :
            select[0:9] == 10'd798 ? table_port[798] :
            select[0:9] == 10'd799 ? table_port[799] :
            select[0:9] == 10'd800 ? table_port[800] :
            select[0:9] == 10'd801 ? table_port[801] :
            select[0:9] == 10'd802 ? table_port[802] :
            select[0:9] == 10'd803 ? table_port[803] :
            select[0:9] == 10'd804 ? table_port[804] :
            select[0:9] == 10'd805 ? table_port[805] :
            select[0:9] == 10'd806 ? table_port[806] :
            select[0:9] == 10'd807 ? table_port[807] :
            select[0:9] == 10'd808 ? table_port[808] :
            select[0:9] == 10'd809 ? table_port[809] :
            select[0:9] == 10'd810 ? table_port[810] :
            select[0:9] == 10'd811 ? table_port[811] :
            select[0:9] == 10'd812 ? table_port[812] :
            select[0:9] == 10'd813 ? table_port[813] :
            select[0:9] == 10'd814 ? table_port[814] :
            select[0:9] == 10'd815 ? table_port[815] :
            select[0:9] == 10'd816 ? table_port[816] :
            select[0:9] == 10'd817 ? table_port[817] :
            select[0:9] == 10'd818 ? table_port[818] :
            select[0:9] == 10'd819 ? table_port[819] :
            select[0:9] == 10'd820 ? table_port[820] :
            select[0:9] == 10'd821 ? table_port[821] :
            select[0:9] == 10'd822 ? table_port[822] :
            select[0:9] == 10'd823 ? table_port[823] :
            select[0:9] == 10'd824 ? table_port[824] :
            select[0:9] == 10'd825 ? table_port[825] :
            select[0:9] == 10'd826 ? table_port[826] :
            select[0:9] == 10'd827 ? table_port[827] :
            select[0:9] == 10'd828 ? table_port[828] :
            select[0:9] == 10'd829 ? table_port[829] :
            select[0:9] == 10'd830 ? table_port[830] :
            select[0:9] == 10'd831 ? table_port[831] :
            select[0:9] == 10'd832 ? table_port[832] :
            select[0:9] == 10'd833 ? table_port[833] :
            select[0:9] == 10'd834 ? table_port[834] :
            select[0:9] == 10'd835 ? table_port[835] :
            select[0:9] == 10'd836 ? table_port[836] :
            select[0:9] == 10'd837 ? table_port[837] :
            select[0:9] == 10'd838 ? table_port[838] :
            select[0:9] == 10'd839 ? table_port[839] :
            select[0:9] == 10'd840 ? table_port[840] :
            select[0:9] == 10'd841 ? table_port[841] :
            select[0:9] == 10'd842 ? table_port[842] :
            select[0:9] == 10'd843 ? table_port[843] :
            select[0:9] == 10'd844 ? table_port[844] :
            select[0:9] == 10'd845 ? table_port[845] :
            select[0:9] == 10'd846 ? table_port[846] :
            select[0:9] == 10'd847 ? table_port[847] :
            select[0:9] == 10'd848 ? table_port[848] :
            select[0:9] == 10'd849 ? table_port[849] :
            select[0:9] == 10'd850 ? table_port[850] :
            select[0:9] == 10'd851 ? table_port[851] :
            select[0:9] == 10'd852 ? table_port[852] :
            select[0:9] == 10'd853 ? table_port[853] :
            select[0:9] == 10'd854 ? table_port[854] :
            select[0:9] == 10'd855 ? table_port[855] :
            select[0:9] == 10'd856 ? table_port[856] :
            select[0:9] == 10'd857 ? table_port[857] :
            select[0:9] == 10'd858 ? table_port[858] :
            select[0:9] == 10'd859 ? table_port[859] :
            select[0:9] == 10'd860 ? table_port[860] :
            select[0:9] == 10'd861 ? table_port[861] :
            select[0:9] == 10'd862 ? table_port[862] :
            select[0:9] == 10'd863 ? table_port[863] :
            select[0:9] == 10'd864 ? table_port[864] :
            select[0:9] == 10'd865 ? table_port[865] :
            select[0:9] == 10'd866 ? table_port[866] :
            select[0:9] == 10'd867 ? table_port[867] :
            select[0:9] == 10'd868 ? table_port[868] :
            select[0:9] == 10'd869 ? table_port[869] :
            select[0:9] == 10'd870 ? table_port[870] :
            select[0:9] == 10'd871 ? table_port[871] :
            select[0:9] == 10'd872 ? table_port[872] :
            select[0:9] == 10'd873 ? table_port[873] :
            select[0:9] == 10'd874 ? table_port[874] :
            select[0:9] == 10'd875 ? table_port[875] :
            select[0:9] == 10'd876 ? table_port[876] :
            select[0:9] == 10'd877 ? table_port[877] :
            select[0:9] == 10'd878 ? table_port[878] :
            select[0:9] == 10'd879 ? table_port[879] :
            select[0:9] == 10'd880 ? table_port[880] :
            select[0:9] == 10'd881 ? table_port[881] :
            select[0:9] == 10'd882 ? table_port[882] :
            select[0:9] == 10'd883 ? table_port[883] :
            select[0:9] == 10'd884 ? table_port[884] :
            select[0:9] == 10'd885 ? table_port[885] :
            select[0:9] == 10'd886 ? table_port[886] :
            select[0:9] == 10'd887 ? table_port[887] :
            select[0:9] == 10'd888 ? table_port[888] :
            select[0:9] == 10'd889 ? table_port[889] :
            select[0:9] == 10'd890 ? table_port[890] :
            select[0:9] == 10'd891 ? table_port[891] :
            select[0:9] == 10'd892 ? table_port[892] :
            select[0:9] == 10'd893 ? table_port[893] :
            select[0:9] == 10'd894 ? table_port[894] :
            select[0:9] == 10'd895 ? table_port[895] :
            select[0:9] == 10'd896 ? table_port[896] :
            select[0:9] == 10'd897 ? table_port[897] :
            select[0:9] == 10'd898 ? table_port[898] :
            select[0:9] == 10'd899 ? table_port[899] :
            select[0:9] == 10'd900 ? table_port[900] :
            select[0:9] == 10'd901 ? table_port[901] :
            select[0:9] == 10'd902 ? table_port[902] :
            select[0:9] == 10'd903 ? table_port[903] :
            select[0:9] == 10'd904 ? table_port[904] :
            select[0:9] == 10'd905 ? table_port[905] :
            select[0:9] == 10'd906 ? table_port[906] :
            select[0:9] == 10'd907 ? table_port[907] :
            select[0:9] == 10'd908 ? table_port[908] :
            select[0:9] == 10'd909 ? table_port[909] :
            select[0:9] == 10'd910 ? table_port[910] :
            select[0:9] == 10'd911 ? table_port[911] :
            select[0:9] == 10'd912 ? table_port[912] :
            select[0:9] == 10'd913 ? table_port[913] :
            select[0:9] == 10'd914 ? table_port[914] :
            select[0:9] == 10'd915 ? table_port[915] :
            select[0:9] == 10'd916 ? table_port[916] :
            select[0:9] == 10'd917 ? table_port[917] :
            select[0:9] == 10'd918 ? table_port[918] :
            select[0:9] == 10'd919 ? table_port[919] :
            select[0:9] == 10'd920 ? table_port[920] :
            select[0:9] == 10'd921 ? table_port[921] :
            select[0:9] == 10'd922 ? table_port[922] :
            select[0:9] == 10'd923 ? table_port[923] :
            select[0:9] == 10'd924 ? table_port[924] :
            select[0:9] == 10'd925 ? table_port[925] :
            select[0:9] == 10'd926 ? table_port[926] :
            select[0:9] == 10'd927 ? table_port[927] :
            select[0:9] == 10'd928 ? table_port[928] :
            select[0:9] == 10'd929 ? table_port[929] :
            select[0:9] == 10'd930 ? table_port[930] :
            select[0:9] == 10'd931 ? table_port[931] :
            select[0:9] == 10'd932 ? table_port[932] :
            select[0:9] == 10'd933 ? table_port[933] :
            select[0:9] == 10'd934 ? table_port[934] :
            select[0:9] == 10'd935 ? table_port[935] :
            select[0:9] == 10'd936 ? table_port[936] :
            select[0:9] == 10'd937 ? table_port[937] :
            select[0:9] == 10'd938 ? table_port[938] :
            select[0:9] == 10'd939 ? table_port[939] :
            select[0:9] == 10'd940 ? table_port[940] :
            select[0:9] == 10'd941 ? table_port[941] :
            select[0:9] == 10'd942 ? table_port[942] :
            select[0:9] == 10'd943 ? table_port[943] :
            select[0:9] == 10'd944 ? table_port[944] :
            select[0:9] == 10'd945 ? table_port[945] :
            select[0:9] == 10'd946 ? table_port[946] :
            select[0:9] == 10'd947 ? table_port[947] :
            select[0:9] == 10'd948 ? table_port[948] :
            select[0:9] == 10'd949 ? table_port[949] :
            select[0:9] == 10'd950 ? table_port[950] :
            select[0:9] == 10'd951 ? table_port[951] :
            select[0:9] == 10'd952 ? table_port[952] :
            select[0:9] == 10'd953 ? table_port[953] :
            select[0:9] == 10'd954 ? table_port[954] :
            select[0:9] == 10'd955 ? table_port[955] :
            select[0:9] == 10'd956 ? table_port[956] :
            select[0:9] == 10'd957 ? table_port[957] :
            select[0:9] == 10'd958 ? table_port[958] :
            select[0:9] == 10'd959 ? table_port[959] :
            select[0:9] == 10'd960 ? table_port[960] :
            select[0:9] == 10'd961 ? table_port[961] :
            select[0:9] == 10'd962 ? table_port[962] :
            select[0:9] == 10'd963 ? table_port[963] :
            select[0:9] == 10'd964 ? table_port[964] :
            select[0:9] == 10'd965 ? table_port[965] :
            select[0:9] == 10'd966 ? table_port[966] :
            select[0:9] == 10'd967 ? table_port[967] :
            select[0:9] == 10'd968 ? table_port[968] :
            select[0:9] == 10'd969 ? table_port[969] :
            select[0:9] == 10'd970 ? table_port[970] :
            select[0:9] == 10'd971 ? table_port[971] :
            select[0:9] == 10'd972 ? table_port[972] :
            select[0:9] == 10'd973 ? table_port[973] :
            select[0:9] == 10'd974 ? table_port[974] :
            select[0:9] == 10'd975 ? table_port[975] :
            select[0:9] == 10'd976 ? table_port[976] :
            select[0:9] == 10'd977 ? table_port[977] :
            select[0:9] == 10'd978 ? table_port[978] :
            select[0:9] == 10'd979 ? table_port[979] :
            select[0:9] == 10'd980 ? table_port[980] :
            select[0:9] == 10'd981 ? table_port[981] :
            select[0:9] == 10'd982 ? table_port[982] :
            select[0:9] == 10'd983 ? table_port[983] :
            select[0:9] == 10'd984 ? table_port[984] :
            select[0:9] == 10'd985 ? table_port[985] :
            select[0:9] == 10'd986 ? table_port[986] :
            select[0:9] == 10'd987 ? table_port[987] :
            select[0:9] == 10'd988 ? table_port[988] :
            select[0:9] == 10'd989 ? table_port[989] :
            select[0:9] == 10'd990 ? table_port[990] :
            select[0:9] == 10'd991 ? table_port[991] :
            select[0:9] == 10'd992 ? table_port[992] :
            select[0:9] == 10'd993 ? table_port[993] :
            select[0:9] == 10'd994 ? table_port[994] :
            select[0:9] == 10'd995 ? table_port[995] :
            select[0:9] == 10'd996 ? table_port[996] :
            select[0:9] == 10'd997 ? table_port[997] :
            select[0:9] == 10'd998 ? table_port[998] : table_port[999]); 

endmodule
